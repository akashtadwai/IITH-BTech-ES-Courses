module splice_demo(a, b, c, d, e, f, x, y);
    input [1:0] a, b, c, d, e, f;
    output [1:0] x = {a[0], a[1]};
    output [11:0] y;
    assign {y[11:4], y[1:0], y[3:2]} = {a, b, -{c, d}, ~{e, f}};
endmodule
