
module tb();



endmodule

