module direct(inp, outp);
    input wire inp;
    output wire outp;
    assign outp = inp;
endmodule
